# ====================================================================
#
#      i2c_freescale.cdl
#
#      eCos Freescale Kinetis and ColdFire+ I2C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Tomas Frydrych
# Contributors:
# Date:           2011-11-20
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_interface CYGINT_IO_FREESCALE_I2C_BUS {
    display      "Number of I2C buses"
}

cdl_package CYGPKG_DEVS_I2C_FREESCALE_I2C {
    display       "Freescale I2C driver"
    parent        CYGPKG_IO_I2C
    requires      CYGPKG_IO_I2C
    requires      CYGPKG_HAL_CORTEXM_KINETIS
    include_dir   cyg/io
    description   "
        This package provides a generic I2C device driver for the on-chip
        I2C modules in Freescale Kinetis and ColdFire+ chips."

    compile       -library=libextras.a i2c_freescale.c

    for { set ::bus 0 } { $::bus < 2 } { incr ::bus } {

        cdl_interface CYGINT_IO_FREESCALE_I2C[set ::bus] {
            display "I2C bus [set ::bus] is present"
        }

        cdl_component CYGHWR_DEVS_FREESCALE_I2C[set ::bus] {
            display       "I2C bus [set ::bus]"
            flavor        bool
            description   "Enable I2C bus [set ::bus]"
            requires      CYGPKG_DEVS_I2C_FREESCALE_I2C
            active_if     CYGINT_IO_FREESCALE_I2C[set ::bus]
            implements    CYGINT_IO_FREESCALE_I2C_BUS
            default_value 0

            cdl_component CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK {
                display       "Default I2C bus frequency"
                flavor        data
                description   "
                    The default frequency setting for I2C[set ::bus].
                    If bit 31 is set then the least significant byte contains
                    pre-calculeted frequency divider register setting.
                    Otherwise other bits contain frequency setpoint in \[Hz\]."

                    requires (CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK > 0 &&            \
                             CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK <= 268435455) ||   \
                             (CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK >= 0x80000000 &&  \
                             CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK <= 0x800000FF)

                default_value 100000

                cdl_option CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK_FIT {
                    display       "Fit"
                    flavor        data
                    legal_values  1 2 3
                    default_value 1
                    description   "
                        For a given clock frequency there are several divider
                        register that fit. This option is hints on which fit to end lookup"
                    }

                cdl_option CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_CLOCK_AGR {
                    display       "Aggressive clocking"
                    flavor        data
                    legal_values  0 1
                    default_value 0
                    description   "
                        If the setpoint bus frequency is not available, then if
                        this option is 1 the closest available frequency is
                        picked even if it overclocks. If 0 the closest available
                        frequency frequency not higher than setpoint is picked."
                }
            }

            cdl_component CYGOPT_DEVS_FREESCALE_I2C[set ::bus]_C2 {
                display        "C2 register options"
                flavor         data
                calculated 0x0 |                                     \
                      CYGOPT_DEVS_FREESCALE_I2C[set ::bus]_C2_HDRS << 5

                cdl_option CYGOPT_DEVS_FREESCALE_I2C[set ::bus]_C2_HDRS {
                    display       "High drive select"
                    flavor        bool
                    no_define
                    default_value 0
                }
            }

            cdl_option CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_FLT {
                display         "Glitch filter"
                flavor          data
                default_value   0
                legal_values    { 0 to 31 }
            }
        }
    }

    cdl_option CYGPKG_DEVS_I2C_FREESCALE_I2C_TRACE {
        display       "I2C trace"
        flavor        bool
        default_value 0
        description   "
            Enable I2C transaction trace. Select to debug the driver."
    }

    cdl_component CYGPKG_DEVS_I2C_FREESCALE_I2C_OPTIONS {
        display      "I2C driver build options"
        flavor        none
        description   "
            Package specific build options including control over
            compiler flags used only in building the Freescale I2C bus driver."

        cdl_option CYGPKG_DEVS_I2C_FREESCALE_I2C_CFLAGS_ADD {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Freescale I2C bus driver. These
                flags are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_I2C_FREESCALE_I2C_CFLAGS_REMOVE {
            display       "Suppressed compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Freescale I2C bus driver. These
                flags are removed from the set of global flags if
                present."
        }
    }
}

# EOF i2c_freescale.cdl
