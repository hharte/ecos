# ====================================================================
#
#      flash_strata_v2.cdl
#
#      FLASH memory - Hardware support for Intel Strata Flash
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:   Andrew Lunn
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_STRATA_V2 {
    display       "Intel StrataFLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    implements    CYGHWR_IO_FLASH_DEVICE

    active_if     CYGINT_DEVS_FLASH_STRATA_V2_REQUIRED

    include_dir   cyg/io

    description   "FLASH memory device support for Intel StrataFlash using
                   the V2 driver API"

    cdl_component CYGOPT_DEVS_FLASH_STRATA_V2_LOCKING {
	display       "Flash device implements locking"
	default_value 1
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        description   "
            This option controls whether the driver will include code
            to allow locking and unlocking of blocks."

        cdl_option CYGNUM_DEVS_FLASH_STRATA_V2_MAX_BLOCKS {
             display       "Maximum number of blocks the driver supports" 
             flavor        data
             default_value 128
             description   "
                 The strata devices do not support unlocking an 
                 individual block. Instead it is necassary to unlock
                 all the blocks in one operation and then lock all those
                 blocks that should be blocked. To do this we need an array
                 containing the current status of the blocks. This controls the 
                 size of that array."
        }       
    }

    cdl_option  CYGOPT_DEV_FLASH_STATE_V2_DUMP_UNKNOWN {
        display       "Dump the identification string for unknown devices"
        default_value 0
        description   "
            This option, when enabled, causes the device driver to 
            dump the identification string when it finds a device it cannot
            identify. Seeing this information is useful for debugging when
            the driver fails to recoginise the device. However in normal 
            operation you probably don't want to see this information 
            because it could acutally be another device some other driver
            in the image can driver."
    }
}

