# ====================================================================
#
#      io_flash.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Gary Thomas
## Copyright (C) 2004 Andrew Lunn
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:   woehler
# Date:           2000-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_FLASH {
    display       "FLASH device drivers"
    include_dir   cyg/io
    doc           ref/flash.html
    description   "
        This option enables drivers for basic I/O services on
        flash devices."
    requires CYGPKG_ISOINFRA
    requires CYGINT_ISO_STRING_STRFUNCS

    compile       flash.c
 
    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>"
        puts $::cdl_header "#ifdef CYGDAT_IO_FLASH_DEVICE_HEADER"
        puts $::cdl_header "# include CYGDAT_IO_FLASH_DEVICE_HEADER"
        puts $::cdl_header "#endif "
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE {
        display       "Hardware FLASH device drivers"
        description   "
            This option enables the hardware device drivers
            for the current platform."
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM {
        display       "Hardware FLASH device drivers are not in RAM"
        flavor        booldata
        description   "
            Use of this interface is deprecated.
            Drivers should make sure that the functions are
            linked to RAM by putting them in .2ram sections."
            requires !CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM
    }

    cdl_interface CYGHWR_IO_FLASH_BLOCK_LOCKING {
        display       "Hardware can support block locking"
        flavor        booldata
        description   "
            This option will be enabled by devices which can support
            locking (write-protection) of individual blocks."
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE_LEGACY {
        display       "Hardware driver uses the legacy interface"
        flavor        booldata
        description   "
            The flash device driver implements the legacy interface to the 
            flash library"
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE_V2 {
        display       "Hardware driver uses the V2 interface"
        flavor        booldata
        description   "
            The flash device driver implements the V2 interface to the 
            flash library"
    }
        
    cdl_option CYGSEM_IO_FLASH_READ_INDIRECT {
        display       "Hardware cannot support direct access to FLASH memory"
        flavor        bool
        default_value 0
        requires      { !CYGSEM_IO_FLASH_VERIFY_PROGRAM }
        description   "
            This option will be asserted by devices which cannot support
            direct access to the FLASH memory contents (e.g. EEPROM or NAND
            devices).  In these cases, the driver must provide an appropriate
            hardware access function."
    }

    cdl_option CYGSEM_IO_FLASH_CHATTER {
        display          "Display status messages during flash operations"
        flavor           bool
        default_value    1
        description      "
           Selecting this option will cause the drivers to print status
           messages as various flash operations are undertaken."
    }

    cdl_option CYGSEM_IO_FLASH_VERIFY_PROGRAM {
        display          "Verify data programmed to flash"
        flavor           bool
        default_value    1
        description      "
           Selecting this option will cause verification of data
           programmed to flash."
    }

    cdl_option CYGSEM_IO_FLASH_SOFT_WRITE_PROTECT {
        display          "Platform has flash soft DIP switch write-protect"
        flavor           bool
        default_value    0
        description      "
           Selecting this option will cause the state of a hardware jumper or
           dipswitch to be read by software to determine whether the flash is
           write-protected or not."
    }


    cdl_option CYGSEM_IO_FLASH_LEGACY_API {
        display          "Provide the legacy user API"
        flavor           bool
        default_value    1
        compile          legacy_api.c
        description      "
            Provide an implementation of the lagacy user API. This is mapped 
            onto the new API via a small layer of code"
    }
        
    cdl_option CYGSEM_IO_FLASH_LEGACY_DEVICE_API {
        display          "Provide the legacy device API"
        flavor           bool
        default_value    CYGHWR_IO_FLASH_DEVICE_LEGACY
        compile          -library=libextras.a legacy_dev.c
        description      "
            Provide an implementation of the legacy device API. This can be 
            used to interface to one legacy device."
    }
    
    cdl_component CYGPKG_IO_FLASH_BLOCK_DEVICE {
        display         "Instantiate in I/O block device API"
        flavor          bool
        active_if       CYGPKG_IO
        default_value   0
        compile         -library=libextras.a flashiodev.c
        description     "
                Provides a block device accessible using the standard I/O
                API ( cyg_io_read() etc. )"

        cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_1 {
            display       "Name of flash device 1 block device"
            flavor        data
            default_value { "\"/dev/flash1\"" }
                
            cdl_interface CYGINT_IO_FLASH_BLOCK_CFG_1 {
                  requires 1 == CYGINT_IO_FLASH_BLOCK_CFG_1
                  no_define
            }

            cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_STATIC_1 {
                  display       "Static configuration via offset"
                  default_value 1
                  implements    CYGINT_IO_FLASH_BLOCK_CFG_1
                  description   "
                        This configures the flash device 1 block device
                        with static offset from the base of the first
                        flash device and length"
                        
                  cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_1 {
                      display         "Start offset from flash base"
                      flavor          data
                      default_value   0x100000
                      description     "
                            This gives the offset from the base of flash 
                            of the first flash device which this block device 
                            corresponds to."
                  }
                  cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_1 {
                      display         "Length"
                      flavor          data
                      default_value   0x100000
                      description     "
                            This gives the length of the region of flash given over
                            to this block device."
                  }
            }
            cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_STATIC_ABSOLUTE_1 {
                  display       "Absolute static configuration"
                  default_value 0
                  implements    CYGINT_IO_FLASH_BLOCK_CFG_1
                  description   "
                        This configures the flash device 1 block device
                        with absolute base address and a length"
                        
                   cdl_option CYGNUM_IO_FLASH_BLOCK_ABSOLUTE_START_1 {
                       display         "Start offset from flash base"
                       flavor          data
                       default_value   0x4000000
                       description     "
                             This gives the absolute address in flash which this
                             block device corresponds to."
                   }
                   cdl_option CYGNUM_IO_FLASH_BLOCK_ABSOLUTE_LENGTH_1 {
                       display         "Length"
                       flavor          data
                       default_value   0x100000
                       description     "
                             This gives the length of the region of flash given over
                             to this block device."
                   }
             }
             cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_FIS_1 {
                    display       "Configuration from FIS"
                    default_value 0
                    implements    CYGINT_IO_FLASH_BLOCK_CFG_1
                    description   "
                          This configures the flash device 1 block device
                          from Redboot FIS"
                                       
                     cdl_component CYGDAT_IO_FLASH_BLOCK_FIS_NAME_1 {
                            display       "Name of FIS entry"
                            flavor        data
                            default_value { "\"jffs2\"" }   
                     }
            }        
        }        
        cdl_component CYGSEM_IO_FLASH_BLOCK_DEVICE_2 {
               display       "Implements a second block device"
               default_value 0

               cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_2 {
               display       "Name of flash device 2 block device"
               flavor        data
               default_value { "\"/dev/flash2\"" }
                
               cdl_interface CYGINT_IO_FLASH_BLOCK_CFG_2 {
                             requires 1 == CYGINT_IO_FLASH_BLOCK_CFG_2
                             no_define
               }

               cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_STATIC_2 {
                      display       "Static configuration via offset"
                      default_value 1
                      implements    CYGINT_IO_FLASH_BLOCK_CFG_2
                      description   "
                            This configures the flash device 2 block device
                            with static offset from the base of the first
                            flash device and length"
                        
                      cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_2 {
                            display         "Start offset from flash base"
                            flavor          data
                            default_value   0x100000
                            description     "
                                  This gives the offset from the base of flash 
                                  of the first flash device which this block device 
                                  corresponds to."
                      }
                      cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_2 {
                            display         "Length"
                            flavor          data
                            default_value   0x100000
                            description     "
                                  This gives the length of the region of flash 
                                  given over to this block device."
                      }       
               }
               cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_STATIC_ABSOLUTE_2 {
                      display       "Absolute static configuration"
                      default_value 0
                      implements    CYGINT_IO_FLASH_BLOCK_CFG_2
                      description   "
                            This configures the flash device 2 block device
                            with absolute base address and a length"
                        
                      cdl_option CYGNUM_IO_FLASH_BLOCK_ABSOLUTE_START_2 {
                            display         "Start offset from flash base"
                            flavor          data
                            default_value   0x4000000
                            description     "
                                  This gives the absolute address in flash which this
                                  block device corresponds to."
                      }
                      cdl_option CYGNUM_IO_FLASH_BLOCK_ABSOLUTE_LENGTH_2 {
                            display         "Length"
                            flavor          data
                            default_value   0x100000
                            description     "
                                  This gives the length of the region of flash 
                                  given over to this block device."
                      }
               }

               cdl_component CYGNUM_IO_FLASH_BLOCK_CFG_FIS_2 {
                      display       "Configuration from FIS"
                      default_value 0
                      implements    CYGINT_IO_FLASH_BLOCK_CFG_2
                      description   "
                            This configures the flash device 2 block device
                            from Redboot FIS"
                                       
                      cdl_component CYGDAT_IO_FLASH_BLOCK_FIS_NAME_2 {
                            display       "Name of FIS entry"
                            flavor        data
                            default_value { "\"jffs2-2\"" }   
                      }
               }        
            }
         }
     }
}